VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO SRAM_4x16_1rw
   CLASS BLOCK ;
   SIZE 33.18 BY 53.06 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  17.08 0.0 17.22 0.42 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  20.16 0.0 20.3 0.42 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  22.68 0.0 22.82 0.42 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  25.76 0.0 25.9 0.42 ;
      END
   END din0[3]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 40.6 0.42 40.74 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  11.76 52.64 11.9 53.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  11.2 52.64 11.34 53.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  11.48 52.64 11.62 53.06 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 4.76 0.42 4.9 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 7.28 0.42 7.42 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.52 0.0 9.66 0.42 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 17.08 33.18 17.22 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 15.68 33.18 15.82 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 15.96 33.18 16.1 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 16.24 33.18 16.38 ;
      END
   END dout0[3]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.96 1.96 31.22 2.66 ;
         LAYER metal4 ;
         RECT  30.52 1.96 31.22 51.1 ;
         LAYER metal3 ;
         RECT  1.96 50.4 31.22 51.1 ;
         LAYER metal4 ;
         RECT  1.96 1.96 2.66 51.1 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.56 51.8 32.62 52.5 ;
         LAYER metal4 ;
         RECT  0.56 0.56 1.26 52.5 ;
         LAYER metal4 ;
         RECT  31.92 0.56 32.62 52.5 ;
         LAYER metal3 ;
         RECT  0.56 0.56 32.62 1.26 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 33.04 52.92 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 33.04 52.92 ;
   LAYER  metal3 ;
      RECT  0.56 40.46 33.04 40.88 ;
      RECT  0.14 5.04 0.56 7.14 ;
      RECT  0.14 7.56 0.56 40.46 ;
      RECT  0.56 16.94 32.62 17.36 ;
      RECT  0.56 17.36 32.62 40.46 ;
      RECT  32.62 17.36 33.04 40.46 ;
      RECT  32.62 16.52 33.04 16.94 ;
      RECT  0.56 1.82 1.82 2.8 ;
      RECT  0.56 2.8 1.82 16.94 ;
      RECT  1.82 2.8 31.36 16.94 ;
      RECT  31.36 1.82 32.62 2.8 ;
      RECT  31.36 2.8 32.62 16.94 ;
      RECT  0.56 40.88 1.82 50.26 ;
      RECT  0.56 50.26 1.82 51.24 ;
      RECT  1.82 40.88 31.36 50.26 ;
      RECT  31.36 40.88 33.04 50.26 ;
      RECT  31.36 50.26 33.04 51.24 ;
      RECT  0.14 40.88 0.42 51.66 ;
      RECT  0.14 51.66 0.42 52.64 ;
      RECT  0.14 52.64 0.42 52.92 ;
      RECT  0.42 40.88 0.56 51.66 ;
      RECT  0.42 52.64 0.56 52.92 ;
      RECT  0.56 51.24 1.82 51.66 ;
      RECT  0.56 52.64 1.82 52.92 ;
      RECT  1.82 51.24 31.36 51.66 ;
      RECT  1.82 52.64 31.36 52.92 ;
      RECT  31.36 51.24 32.76 51.66 ;
      RECT  31.36 52.64 32.76 52.92 ;
      RECT  32.76 51.24 33.04 51.66 ;
      RECT  32.76 51.66 33.04 52.64 ;
      RECT  32.76 52.64 33.04 52.92 ;
      RECT  0.14 0.14 0.42 0.42 ;
      RECT  0.14 0.42 0.42 1.4 ;
      RECT  0.14 1.4 0.42 4.62 ;
      RECT  0.42 0.14 0.56 0.42 ;
      RECT  0.42 1.4 0.56 4.62 ;
      RECT  32.62 0.14 32.76 0.42 ;
      RECT  32.62 1.4 32.76 15.54 ;
      RECT  32.76 0.14 33.04 0.42 ;
      RECT  32.76 0.42 33.04 1.4 ;
      RECT  32.76 1.4 33.04 15.54 ;
      RECT  0.56 0.14 1.82 0.42 ;
      RECT  0.56 1.4 1.82 1.82 ;
      RECT  1.82 0.14 31.36 0.42 ;
      RECT  1.82 1.4 31.36 1.82 ;
      RECT  31.36 0.14 32.62 0.42 ;
      RECT  31.36 1.4 32.62 1.82 ;
   LAYER  metal4 ;
      RECT  16.8 0.7 17.5 52.92 ;
      RECT  17.5 0.14 19.88 0.7 ;
      RECT  20.58 0.14 22.4 0.7 ;
      RECT  23.1 0.14 25.48 0.7 ;
      RECT  11.48 0.7 12.18 52.36 ;
      RECT  12.18 0.7 16.8 52.36 ;
      RECT  12.18 52.36 16.8 52.92 ;
      RECT  9.94 0.14 16.8 0.7 ;
      RECT  17.5 0.7 30.24 1.68 ;
      RECT  17.5 1.68 30.24 51.38 ;
      RECT  17.5 51.38 30.24 52.92 ;
      RECT  30.24 0.7 31.5 1.68 ;
      RECT  30.24 51.38 31.5 52.92 ;
      RECT  1.68 0.7 2.94 1.68 ;
      RECT  1.68 51.38 2.94 52.36 ;
      RECT  2.94 0.7 11.48 1.68 ;
      RECT  2.94 1.68 11.48 51.38 ;
      RECT  2.94 51.38 11.48 52.36 ;
      RECT  0.14 52.36 0.28 52.78 ;
      RECT  0.14 52.78 0.28 52.92 ;
      RECT  0.28 52.78 1.54 52.92 ;
      RECT  1.54 52.36 10.92 52.78 ;
      RECT  1.54 52.78 10.92 52.92 ;
      RECT  0.14 0.14 0.28 0.28 ;
      RECT  0.14 0.28 0.28 0.7 ;
      RECT  0.28 0.14 1.54 0.28 ;
      RECT  1.54 0.14 9.24 0.28 ;
      RECT  1.54 0.28 9.24 0.7 ;
      RECT  0.14 0.7 0.28 1.68 ;
      RECT  1.54 0.7 1.68 1.68 ;
      RECT  0.14 1.68 0.28 51.38 ;
      RECT  1.54 1.68 1.68 51.38 ;
      RECT  0.14 51.38 0.28 52.36 ;
      RECT  1.54 51.38 1.68 52.36 ;
      RECT  26.18 0.14 31.64 0.28 ;
      RECT  26.18 0.28 31.64 0.7 ;
      RECT  31.64 0.14 32.9 0.28 ;
      RECT  32.9 0.14 33.04 0.28 ;
      RECT  32.9 0.28 33.04 0.7 ;
      RECT  31.5 0.7 31.64 1.68 ;
      RECT  32.9 0.7 33.04 1.68 ;
      RECT  31.5 1.68 31.64 51.38 ;
      RECT  32.9 1.68 33.04 51.38 ;
      RECT  31.5 51.38 31.64 52.78 ;
      RECT  31.5 52.78 31.64 52.92 ;
      RECT  31.64 52.78 32.9 52.92 ;
      RECT  32.9 51.38 33.04 52.78 ;
      RECT  32.9 52.78 33.04 52.92 ;
   END
END    SRAM_4x16_1rw
END    LIBRARY
