VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO SRAM_2x32_1rw
   CLASS BLOCK ;
   SIZE 33.18 BY 52.78 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  20.16 0.0 20.3 0.42 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  22.68 0.0 22.82 0.42 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  17.36 0.0 17.5 0.42 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 40.6 0.42 40.74 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  10.92 52.36 11.06 52.78 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  11.2 52.36 11.34 52.78 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  11.48 52.36 11.62 52.78 ;
      END
   END addr0[4]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 4.2 0.42 4.34 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 7.0 0.42 7.14 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  9.8 0.0 9.94 0.42 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 12.88 33.18 13.02 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  32.76 13.16 33.18 13.3 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.96 1.96 31.22 2.66 ;
         LAYER metal4 ;
         RECT  30.52 1.96 31.22 50.82 ;
         LAYER metal3 ;
         RECT  1.96 50.12 31.22 50.82 ;
         LAYER metal4 ;
         RECT  1.96 1.96 2.66 50.82 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  31.92 0.56 32.62 52.22 ;
         LAYER metal3 ;
         RECT  0.56 51.52 32.62 52.22 ;
         LAYER metal4 ;
         RECT  0.56 0.56 1.26 52.22 ;
         LAYER metal3 ;
         RECT  0.56 0.56 32.62 1.26 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 33.04 52.64 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 33.04 52.64 ;
   LAYER  metal3 ;
      RECT  0.56 40.46 33.04 40.88 ;
      RECT  0.14 4.48 0.56 6.86 ;
      RECT  0.14 7.28 0.56 40.46 ;
      RECT  0.56 12.74 32.62 13.16 ;
      RECT  0.56 13.16 32.62 40.46 ;
      RECT  32.62 13.44 33.04 40.46 ;
      RECT  0.56 1.82 1.82 2.8 ;
      RECT  0.56 2.8 1.82 12.74 ;
      RECT  1.82 2.8 31.36 12.74 ;
      RECT  31.36 1.82 32.62 2.8 ;
      RECT  31.36 2.8 32.62 12.74 ;
      RECT  0.56 40.88 1.82 49.98 ;
      RECT  0.56 49.98 1.82 50.96 ;
      RECT  1.82 40.88 31.36 49.98 ;
      RECT  31.36 40.88 33.04 49.98 ;
      RECT  31.36 49.98 33.04 50.96 ;
      RECT  0.14 40.88 0.42 51.38 ;
      RECT  0.14 51.38 0.42 52.36 ;
      RECT  0.14 52.36 0.42 52.64 ;
      RECT  0.42 40.88 0.56 51.38 ;
      RECT  0.42 52.36 0.56 52.64 ;
      RECT  0.56 50.96 1.82 51.38 ;
      RECT  0.56 52.36 1.82 52.64 ;
      RECT  1.82 50.96 31.36 51.38 ;
      RECT  1.82 52.36 31.36 52.64 ;
      RECT  31.36 50.96 32.76 51.38 ;
      RECT  31.36 52.36 32.76 52.64 ;
      RECT  32.76 50.96 33.04 51.38 ;
      RECT  32.76 51.38 33.04 52.36 ;
      RECT  32.76 52.36 33.04 52.64 ;
      RECT  0.14 0.14 0.42 0.42 ;
      RECT  0.14 0.42 0.42 1.4 ;
      RECT  0.14 1.4 0.42 4.06 ;
      RECT  0.42 0.14 0.56 0.42 ;
      RECT  0.42 1.4 0.56 4.06 ;
      RECT  32.62 0.14 32.76 0.42 ;
      RECT  32.62 1.4 32.76 12.74 ;
      RECT  32.76 0.14 33.04 0.42 ;
      RECT  32.76 0.42 33.04 1.4 ;
      RECT  32.76 1.4 33.04 12.74 ;
      RECT  0.56 0.14 1.82 0.42 ;
      RECT  0.56 1.4 1.82 1.82 ;
      RECT  1.82 0.14 31.36 0.42 ;
      RECT  1.82 1.4 31.36 1.82 ;
      RECT  31.36 0.14 32.62 0.42 ;
      RECT  31.36 1.4 32.62 1.82 ;
   LAYER  metal4 ;
      RECT  19.88 0.7 20.58 52.64 ;
      RECT  20.58 0.14 22.4 0.7 ;
      RECT  17.78 0.14 19.88 0.7 ;
      RECT  10.64 0.7 11.34 52.08 ;
      RECT  11.34 0.7 19.88 52.08 ;
      RECT  11.9 52.08 19.88 52.64 ;
      RECT  10.22 0.14 17.08 0.7 ;
      RECT  20.58 0.7 30.24 1.68 ;
      RECT  20.58 1.68 30.24 51.1 ;
      RECT  20.58 51.1 30.24 52.64 ;
      RECT  30.24 0.7 31.5 1.68 ;
      RECT  30.24 51.1 31.5 52.64 ;
      RECT  1.68 0.7 2.94 1.68 ;
      RECT  1.68 51.1 2.94 52.08 ;
      RECT  2.94 0.7 10.64 1.68 ;
      RECT  2.94 1.68 10.64 51.1 ;
      RECT  2.94 51.1 10.64 52.08 ;
      RECT  23.1 0.14 31.64 0.28 ;
      RECT  23.1 0.28 31.64 0.7 ;
      RECT  31.64 0.14 32.9 0.28 ;
      RECT  32.9 0.14 33.04 0.28 ;
      RECT  32.9 0.28 33.04 0.7 ;
      RECT  31.5 0.7 31.64 1.68 ;
      RECT  32.9 0.7 33.04 1.68 ;
      RECT  31.5 1.68 31.64 51.1 ;
      RECT  32.9 1.68 33.04 51.1 ;
      RECT  31.5 51.1 31.64 52.5 ;
      RECT  31.5 52.5 31.64 52.64 ;
      RECT  31.64 52.5 32.9 52.64 ;
      RECT  32.9 51.1 33.04 52.5 ;
      RECT  32.9 52.5 33.04 52.64 ;
      RECT  0.14 52.08 0.28 52.5 ;
      RECT  0.14 52.5 0.28 52.64 ;
      RECT  0.28 52.5 1.54 52.64 ;
      RECT  1.54 52.08 10.64 52.5 ;
      RECT  1.54 52.5 10.64 52.64 ;
      RECT  0.14 0.14 0.28 0.28 ;
      RECT  0.14 0.28 0.28 0.7 ;
      RECT  0.28 0.14 1.54 0.28 ;
      RECT  1.54 0.14 9.52 0.28 ;
      RECT  1.54 0.28 9.52 0.7 ;
      RECT  0.14 0.7 0.28 1.68 ;
      RECT  1.54 0.7 1.68 1.68 ;
      RECT  0.14 1.68 0.28 51.1 ;
      RECT  1.54 1.68 1.68 51.1 ;
      RECT  0.14 51.1 0.28 52.08 ;
      RECT  1.54 51.1 1.68 52.08 ;
   END
END    SRAM_2x32_1rw
END    LIBRARY
